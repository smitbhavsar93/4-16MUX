library verilog;
use verilog.vl_types.all;
entity dec4to16_vlg_vec_tst is
end dec4to16_vlg_vec_tst;
